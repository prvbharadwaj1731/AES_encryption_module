module MixColumns(
    input [7:0] data_in [3:0][3:0],
    output [7:0] data_out [3:0][3:0]
    );
    



endmodule


//----------------------------------------------------------------------------------------------


